module IFID(
    instr_i,
    instr_o
);

input [31:0] instr_i;
output [31:0] instr_o;


assign instr_o = instr_i;

endmodule
